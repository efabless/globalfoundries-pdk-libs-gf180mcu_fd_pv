
* cell sample_pfet_06v0_dn
.SUBCKT sample_pfet_06v0_dn
* net 1 I1_default_G
* net 2 I1_default_S
* net 3 gnd!
* net 4 I1_default_D
* net 5 I1_lin_default_tapCntRows_4_R0_G
* net 6 I1_lin_default_tapCntRows_0_R0_G
* net 7 I1_lin_default_tapCntRows_1_R0_G
* net 8 I1_lin_default_tapCntRows_2_R0_G
* net 9 I1_lin_default_tapCntRows_3_R0_G
* net 10 I1_lin_default_tapCntRows_0_R0_S
* net 11 I1_lin_default_tapCntRows_4_R0_D
* net 12 I1_lin_default_tapCntRows_0_R0_D
* net 13 I1_lin_default_tapCntRows_1_R0_S
* net 14 I1_lin_default_tapCntRows_4_R0_S
* net 15 I1_lin_default_tapCntRows_3_R0_D
* net 16 I1_lin_default_tapCntRows_1_R0_D
* net 17 I1_lin_default_tapCntRows_2_R0_S
* net 18 I1_lin_default_tapCntRows_2_R0_D
* net 19 I1_lin_default_tapCntRows_3_R0_S
* net 20 I1_lin_default_bottomTap_0_R0_G
* net 21 I1_lin_default_bottomTap_0_R0_S
* net 22 I1_lin_default_bottomTap_0_R0_D
* net 23 I1_lin_default_topTap_0_R0_G
* net 24 I1_lin_default_topTap_0_R0_D
* net 25 I1_lin_default_topTap_0_R0_S
* net 26 I1_lin_default_rightTap_0_R0_G
* net 27 I1_lin_default_rightTap_0_R0_S
* net 28 I1_lin_default_rightTap_0_R0_D
* net 29 I1_lin_default_leftTap_0_R0_S
* net 30 I1_lin_default_leftTap_0_R0_D
* net 31 I1_lin_default_leftTap_0_R0_G
* net 32 I1_lin_default_bodytie_1_R0_G
* net 33 I1_lin_default_bodytie_0_R0_G
* net 34 I1_lin_default_bodytie_0_R0_S
* net 35 I1_lin_default_bodytie_0_R0_D
* net 36 I1_lin_default_bodytie_1_R0_D
* net 37 I1_lin_default_bodytie_1_R0_S
* net 38 I1_lin_default_sdConn_0_R0_G
* net 39 I1_lin_default_sdConn_1_R0_G
* net 40 I1_lin_default_sdConn_2_R0_G
* net 41 I1_lin_default_sdWidth_9_R0_G
* net 42 I1_lin_default_sdConn_0_R0_S
* net 43 I1_lin_default_sdConn_0_R0_D
* net 44 I1_lin_default_sdConn_1_R0_S
* net 45 I1_lin_default_sdConn_2_R0_D
* net 46 I1_lin_default_sdConn_1_R0_D
* net 47 I1_lin_default_sdConn_2_R0_S
* net 48 I1_lin_default_sdWidth_0_R0_G
* net 49 I1_lin_default_sdWidth_1_R0_G
* net 50 I1_lin_default_sdWidth_2_R0_G
* net 51 I1_lin_default_sdWidth_3_R0_G
* net 52 I1_lin_default_sdWidth_4_R0_G
* net 53 I1_lin_default_sdWidth_5_R0_G
* net 54 I1_lin_default_sdWidth_6_R0_G
* net 55 I1_lin_default_sdWidth_7_R0_G
* net 56 I1_lin_default_sdWidth_8_R0_G
* net 57 I1_lin_default_sdWidth_0_R0_S
* net 58 I1_lin_default_sdWidth_1_R0_S
* net 59 I1_lin_default_sdWidth_0_R0_D
* net 60 I1_lin_default_sdWidth_2_R0_S
* net 61 I1_lin_default_sdWidth_9_R0_D
* net 62 I1_lin_default_sdWidth_1_R0_D
* net 63 I1_lin_default_gateConn_2_R0_G
* net 64 I1_lin_default_sdWidth_3_R0_S
* net 65 I1_lin_default_sdWidth_2_R0_D
* net 66 I1_lin_default_sdWidth_4_R0_S
* net 67 I1_lin_default_sdWidth_3_R0_D
* net 68 I1_lin_default_sdWidth_5_R0_S
* net 69 I1_lin_default_sdWidth_4_R0_D
* net 70 I1_lin_default_sdWidth_6_R0_S
* net 71 I1_lin_default_sdWidth_5_R0_D
* net 72 I1_lin_default_sdWidth_7_R0_S
* net 73 I1_lin_default_sdWidth_6_R0_D
* net 74 I1_lin_default_sdWidth_8_R0_S
* net 75 I1_lin_default_sdWidth_7_R0_D
* net 76 I1_lin_default_sdWidth_9_R0_S
* net 77 I1_lin_default_sdWidth_8_R0_D
* net 78 I1_lin_default_gateConn_1_R0_G
* net 79 I1_lin_default_gateConn_0_R0_G
* net 80 I1_lin_default_gateConn_0_R0_S
* net 81 I1_lin_default_gateConn_2_R0_S
* net 82 I1_lin_default_gateConn_1_R0_S
* net 83 I1_lin_default_gateConn_0_R0_D
* net 84 I1_lin_default_gateConn_2_R0_D
* net 85 I1_lin_default_gateConn_1_R0_D
* net 86 I1_lin_default_calculatedParam_0_R0_G
* net 87 I1_lin_default_calculatedParam_1_R0_G
* net 88 I1_lin_default_calculatedParam_2_R0_G
* net 89 I1_lin_default_calculatedParam_2_R0_D
* net 90 I1_lin_default_calculatedParam_0_R0_S
* net 91 I1_lin_default_calculatedParam_1_R0_S
* net 92 I1_lin_default_calculatedParam_0_R0_D
* net 93 I1_lin_default_calculatedParam_2_R0_S
* net 94 I1_lin_default_calculatedParam_1_R0_D
* net 95 I1_lin_default_m_1_R0_G
* net 96 I1_lin_default_m_2_R0_G
* net 97 I1_lin_default_m_0_R0_G
* net 98 I1_lin_default_m_0_R0_S
* net 99 I1_lin_default_m_1_R0_S
* net 100 I1_lin_default_m_0_R0_D
* net 101 I1_lin_default_m_2_R0_S
* net 102 I1_lin_default_m_1_R0_D
* net 103 I1_lin_default_m_2_R0_D
* net 104 I1_lin_default_nf_0_R0_G
* net 105 I1_lin_default_nf_1_R0_G
* net 106 I1_lin_default_nf_2_R0_G
* net 107 I1_lin_default_nf_0_R0_S
* net 108 I1_lin_default_nf_0_R0_D
* net 109 I1_lin_default_nf_2_R0_D
* net 110 I1_lin_default_nf_1_R0_S
* net 111 I1_lin_default_nf_2_R0_S
* net 112 I1_lin_default_nf_1_R0_D
* net 113 I1_lin_default_l_0_R0_G
* net 114 I1_lin_default_l_1_R0_G
* net 115 I1_lin_default_l_2_R0_G
* net 116 I1_lin_default_l_3_R0_G
* net 117 I1_lin_default_l_4_R0_G
* net 118 I1_lin_default_l_5_R0_G
* net 119 I1_lin_default_l_6_R0_G
* net 120 I1_lin_default_l_7_R0_G
* net 121 I1_lin_default_l_8_R0_G
* net 122 I1_lin_default_l_9_R0_G
* net 123 I1_lin_default_l_10_R0_G
* net 124 I1_lin_default_l_11_R0_G
* net 125 I1_lin_default_l_12_R0_G
* net 126 I1_lin_default_l_13_R0_G
* net 127 I1_lin_default_l_14_R0_G
* net 128 I1_lin_default_l_15_R0_G
* net 129 I1_lin_default_l_16_R0_G
* net 130 I1_lin_default_l_17_R0_G
* net 131 I1_lin_default_l_18_R0_G
* net 132 I1_lin_default_l_19_R0_G
* net 133 I1_lin_default_l_20_R0_G
* net 134 I1_lin_default_l_21_R0_G
* net 135 I1_lin_default_l_22_R0_G
* net 136 I1_lin_default_l_23_R0_G
* net 137 I1_lin_default_l_24_R0_G
* net 138 I1_lin_default_l_25_R0_G
* net 139 I1_lin_default_l_0_R0_S
* net 140 I1_lin_default_l_25_R0_D
* net 141 I1_lin_default_l_0_R0_D
* net 142 I1_lin_default_l_1_R0_S
* net 143 I1_lin_default_l_2_R0_S
* net 144 I1_lin_default_l_1_R0_D
* net 145 I1_lin_default_l_3_R0_S
* net 146 I1_lin_default_l_2_R0_D
* net 147 I1_lin_default_l_4_R0_S
* net 148 I1_lin_default_l_3_R0_D
* net 149 I1_lin_default_l_5_R0_S
* net 150 I1_lin_default_l_4_R0_D
* net 151 I1_lin_default_l_6_R0_S
* net 152 I1_lin_default_l_5_R0_D
* net 153 I1_lin_default_l_7_R0_S
* net 154 I1_lin_default_l_6_R0_D
* net 155 I1_lin_default_l_8_R0_S
* net 156 I1_lin_default_l_7_R0_D
* net 157 I1_lin_default_l_9_R0_S
* net 158 I1_lin_default_l_8_R0_D
* net 159 I1_lin_default_l_10_R0_S
* net 160 I1_lin_default_l_9_R0_D
* net 161 I1_lin_default_l_11_R0_S
* net 162 I1_lin_default_l_10_R0_D
* net 163 I1_lin_default_l_12_R0_S
* net 164 I1_lin_default_l_11_R0_D
* net 165 I1_lin_default_l_13_R0_S
* net 166 I1_lin_default_l_12_R0_D
* net 167 I1_lin_default_l_14_R0_S
* net 168 I1_lin_default_l_13_R0_D
* net 169 I1_lin_default_l_15_R0_S
* net 170 I1_lin_default_l_14_R0_D
* net 171 I1_lin_default_l_16_R0_S
* net 172 I1_lin_default_l_15_R0_D
* net 173 I1_lin_default_l_17_R0_S
* net 174 I1_lin_default_l_16_R0_D
* net 175 I1_lin_default_l_18_R0_S
* net 176 I1_lin_default_l_17_R0_D
* net 177 I1_lin_default_l_19_R0_S
* net 178 I1_lin_default_l_18_R0_D
* net 179 I1_lin_default_l_20_R0_S
* net 180 I1_lin_default_l_19_R0_D
* net 181 I1_lin_default_l_21_R0_S
* net 182 I1_lin_default_l_20_R0_D
* net 183 I1_lin_default_l_22_R0_S
* net 184 I1_lin_default_l_21_R0_D
* net 185 I1_lin_default_l_23_R0_S
* net 186 I1_lin_default_l_22_R0_D
* net 187 I1_lin_default_l_24_R0_S
* net 188 I1_lin_default_l_23_R0_D
* net 189 I1_lin_default_l_25_R0_S
* net 190 I1_lin_default_l_24_R0_D
* net 191 I1_lin_default_fingerW_0_R0_D
* net 192 I1_lin_default_fingerW_0_R0_S
* net 193 I1_lin_default_fingerW_0_R0_G
* net 194 I1_lin_default_fingerW_1_R0_G
* net 195 I1_lin_default_fingerW_2_R0_G
* net 196 I1_lin_default_fingerW_3_R0_G
* net 197 I1_lin_default_fingerW_4_R0_G
* net 198 I1_lin_default_fingerW_5_R0_G
* net 199 I1_lin_default_fingerW_6_R0_G
* net 200 I1_lin_default_fingerW_7_R0_G
* net 201 I1_lin_default_fingerW_8_R0_G
* net 202 I1_lin_default_fingerW_9_R0_G
* net 203 I1_lin_default_fingerW_10_R0_G
* net 204 I1_lin_default_fingerW_11_R0_G
* net 205 I1_lin_default_fingerW_12_R0_G
* net 206 I1_lin_default_fingerW_13_R0_G
* net 207 I1_lin_default_fingerW_14_R0_G
* net 208 I1_lin_default_fingerW_15_R0_G
* net 209 I1_lin_default_fingerW_16_R0_G
* net 210 I1_lin_default_fingerW_17_R0_G
* net 211 I1_lin_default_fingerW_18_R0_G
* net 212 I1_lin_default_fingerW_19_R0_G
* net 213 I1_lin_default_fingerW_20_R0_G
* net 214 I1_lin_default_fingerW_21_R0_G
* net 215 I1_lin_default_fingerW_22_R0_G
* net 216 I1_lin_default_fingerW_23_R0_G
* net 217 I1_lin_default_fingerW_24_R0_G
* net 218 I1_lin_default_fingerW_25_R0_G
* net 219 I1_lin_default_fingerW_26_R0_G
* net 220 I1_lin_default_fingerW_27_R0_G
* net 221 I1_lin_default_fingerW_28_R0_G
* net 222 I1_lin_default_fingerW_29_R0_G
* net 223 I1_lin_default_fingerW_30_R0_G
* net 224 I1_lin_default_fingerW_31_R0_G
* net 225 I1_lin_default_fingerW_1_R0_S
* net 226 I1_lin_default_fingerW_2_R0_S
* net 227 I1_lin_default_fingerW_1_R0_D
* net 228 I1_lin_default_fingerW_3_R0_S
* net 229 I1_lin_default_fingerW_2_R0_D
* net 230 I1_lin_default_fingerW_4_R0_S
* net 231 I1_lin_default_fingerW_3_R0_D
* net 232 I1_lin_default_fingerW_5_R0_S
* net 233 I1_lin_default_fingerW_4_R0_D
* net 234 I1_lin_default_fingerW_6_R0_S
* net 235 I1_lin_default_fingerW_5_R0_D
* net 236 I1_lin_default_fingerW_7_R0_S
* net 237 I1_lin_default_fingerW_6_R0_D
* net 238 I1_lin_default_fingerW_8_R0_S
* net 239 I1_lin_default_fingerW_7_R0_D
* net 240 I1_lin_default_fingerW_9_R0_S
* net 241 I1_lin_default_fingerW_8_R0_D
* net 242 I1_lin_default_fingerW_10_R0_S
* net 243 I1_lin_default_fingerW_9_R0_D
* net 244 I1_lin_default_fingerW_11_R0_S
* net 245 I1_lin_default_fingerW_10_R0_D
* net 246 I1_lin_default_fingerW_12_R0_S
* net 247 I1_lin_default_fingerW_11_R0_D
* net 248 I1_lin_default_fingerW_13_R0_S
* net 249 I1_lin_default_fingerW_12_R0_D
* net 250 I1_lin_default_fingerW_14_R0_S
* net 251 I1_lin_default_fingerW_13_R0_D
* net 252 I1_lin_default_fingerW_15_R0_S
* net 253 I1_lin_default_fingerW_14_R0_D
* net 254 I1_lin_default_fingerW_16_R0_S
* net 255 I1_lin_default_fingerW_15_R0_D
* net 256 I1_lin_default_fingerW_17_R0_S
* net 257 I1_lin_default_fingerW_16_R0_D
* net 258 I1_lin_default_fingerW_18_R0_S
* net 259 I1_lin_default_fingerW_17_R0_D
* net 260 I1_lin_default_fingerW_19_R0_S
* net 261 I1_lin_default_fingerW_18_R0_D
* net 262 I1_lin_default_fingerW_20_R0_S
* net 263 I1_lin_default_fingerW_19_R0_D
* net 264 I1_lin_default_fingerW_21_R0_S
* net 265 I1_lin_default_fingerW_20_R0_D
* net 266 I1_lin_default_fingerW_22_R0_S
* net 267 I1_lin_default_fingerW_21_R0_D
* net 268 I1_lin_default_fingerW_23_R0_S
* net 269 I1_lin_default_fingerW_22_R0_D
* net 270 I1_lin_default_fingerW_24_R0_S
* net 271 I1_lin_default_fingerW_23_R0_D
* net 272 I1_lin_default_fingerW_25_R0_S
* net 273 I1_lin_default_fingerW_24_R0_D
* net 274 I1_lin_default_fingerW_26_R0_S
* net 275 I1_lin_default_fingerW_25_R0_D
* net 276 I1_lin_default_fingerW_27_R0_S
* net 277 I1_lin_default_fingerW_26_R0_D
* net 278 I1_lin_default_fingerW_28_R0_S
* net 279 I1_lin_default_fingerW_27_R0_D
* net 280 I1_lin_default_fingerW_29_R0_S
* net 281 I1_lin_default_fingerW_28_R0_D
* net 282 I1_lin_default_fingerW_30_R0_S
* net 283 I1_lin_default_fingerW_29_R0_D
* net 284 I1_lin_default_fingerW_31_R0_S
* net 285 I1_lin_default_fingerW_30_R0_D
* net 286 I1_lin_default_fingerW_32_R0_S
* net 287 I1_lin_default_fingerW_31_R0_D
* net 288 I1_lin_default_fingerW_32_R0_D
* net 289 I1_lin_default_fingerW_32_R0_G
* cell instance $1 r0 *1 2.2,1.6
X$1 4 2 1 3 pfet_06v0_dn_CDNS_631264496070
* cell instance $2 r0 *1 9.82,1.92
X$2 3 M1_NACTIVE_CDNS_631264496070
* cell instance $3 r0 *1 40.6,10.2
X$3 3 11 14 5 pfet_06v0_dn_CDNS_6312644960789
* cell instance $4 r0 *1 11.8,10.2
X$4 3 16 13 7 pfet_06v0_dn_CDNS_6312644960788
* cell instance $5 r0 *1 21.4,10.2
X$5 3 18 17 8 pfet_06v0_dn_CDNS_631264496071
* cell instance $6 r0 *1 31,10.2
X$6 3 19 15 9 pfet_06v0_dn_CDNS_631264496072
* cell instance $7 r0 *1 2.2,10.2
X$7 3 12 10 6 pfet_06v0_dn_CDNS_6312644960727
* cell instance $8 r0 *1 2.2,44.6
X$8 3 30 29 31 pfet_06v0_dn_CDNS_631264496077
* cell instance $9 r0 *1 2.2,18.8
X$9 3 22 21 20 pfet_06v0_dn_CDNS_631264496074
* cell instance $10 r0 *1 2.2,27.4
X$10 3 24 25 23 pfet_06v0_dn_CDNS_631264496075
* cell instance $11 r0 *1 2.2,36
X$11 3 28 27 26 pfet_06v0_dn_CDNS_631264496076
* cell instance $12 r0 *1 2.2,53.2
X$12 3 35 34 33 pfet_06v0_dn_CDNS_631264496078
* cell instance $13 r0 *1 11.8,53.2
X$13 3 36 37 32 pfet_06v0_dn_CDNS_631264496073
* cell instance $14 r0 *1 2.2,61.8
X$14 42 43 38 3 pfet_06v0_dn_CDNS_6312644960713
* cell instance $15 r0 *1 21.4,61.8
X$15 47 45 40 3 pfet_06v0_dn_CDNS_6312644960712
* cell instance $16 r0 *1 2.2,70.4
X$16 59 57 48 3 pfet_06v0_dn_CDNS_6312644960715
* cell instance $17 r0 *1 11.8,70.4
X$17 62 58 49 3 pfet_06v0_dn_CDNS_6312644960716
* cell instance $18 r0 *1 21.6,70.4
X$18 65 60 50 3 pfet_06v0_dn_CDNS_6312644960717
* cell instance $19 r0 *1 31.4,70.4
X$19 67 64 51 3 pfet_06v0_dn_CDNS_6312644960718
* cell instance $20 r0 *1 41.6,70.4
X$20 69 66 52 3 pfet_06v0_dn_CDNS_6312644960719
* cell instance $21 r0 *1 51.8,70.4
X$21 71 68 53 3 pfet_06v0_dn_CDNS_6312644960720
* cell instance $22 r0 *1 62.2,70.4
X$22 73 70 54 3 pfet_06v0_dn_CDNS_6312644960721
* cell instance $23 r0 *1 72.8,70.4
X$23 75 72 55 3 pfet_06v0_dn_CDNS_6312644960722
* cell instance $24 r0 *1 83.8,70.4
X$24 77 74 56 3 pfet_06v0_dn_CDNS_6312644960723
* cell instance $25 r0 *1 95,70.4
X$25 61 76 41 3 pfet_06v0_dn_CDNS_6312644960711
* cell instance $26 r0 *1 2.2,79
X$26 83 80 79 3 pfet_06v0_dn_CDNS_6312644960714
* cell instance $27 r0 *1 11.8,87.6
X$27 91 94 87 3 pfet_06v0_dn_CDNS_6312644960726
* cell instance $28 r0 *1 11.8,79
X$28 85 82 78 3 pfet_06v0_dn_CDNS_6312644960725
* cell instance $29 r0 *1 21.4,79
X$29 63 84 81 3 pfet_06v0_dn_CDNS_6312644960724
* cell instance $30 r0 *1 31.81,87.6
X$30 93 89 88 3 pfet_06v0_dn_CDNS_6312644960790
* cell instance $31 r0 *1 -25.015,96.2
X$31 102 99 95 3 pfet_06v0_dn_CDNS_631264496079
* cell instance $32 r0 *1 -15.415,96.2
X$32 101 103 96 3 pfet_06v0_dn_CDNS_6312644960728
* cell instance $33 r0 *1 11.8,104.8
X$33 112 110 105 3 pfet_06v0_dn_CDNS_6312644960729
* cell instance $34 r0 *1 74.8,104.8
X$34 109 111 106 3 pfet_06v0_dn_CDNS_6312644960710
* cell instance $35 r0 *1 2.2,113.4
X$35 141 139 113 3 pfet_06v0_dn_CDNS_6312644960730
* cell instance $36 r0 *1 11.8,113.4
X$36 144 142 114 3 pfet_06v0_dn_CDNS_6312644960731
* cell instance $37 r0 *1 21.6,113.4
X$37 146 143 115 3 pfet_06v0_dn_CDNS_6312644960732
* cell instance $38 r0 *1 31.4,113.4
X$38 148 145 116 3 pfet_06v0_dn_CDNS_6312644960733
* cell instance $39 r0 *1 41.4,113.4
X$39 150 147 117 3 pfet_06v0_dn_CDNS_6312644960734
* cell instance $40 r0 *1 51.6,113.4
X$40 152 149 118 3 pfet_06v0_dn_CDNS_6312644960735
* cell instance $41 r0 *1 62,113.4
X$41 154 151 119 3 pfet_06v0_dn_CDNS_6312644960736
* cell instance $42 r0 *1 72.8,113.4
X$42 156 153 120 3 pfet_06v0_dn_CDNS_6312644960737
* cell instance $43 r0 *1 83.8,113.4
X$43 158 155 121 3 pfet_06v0_dn_CDNS_6312644960738
* cell instance $44 r0 *1 95.2,113.4
X$44 160 157 122 3 pfet_06v0_dn_CDNS_6312644960739
* cell instance $45 r0 *1 107.2,113.4
X$45 162 159 123 3 pfet_06v0_dn_CDNS_6312644960740
* cell instance $46 r0 *1 119.6,113.4
X$46 164 161 124 3 pfet_06v0_dn_CDNS_6312644960741
* cell instance $47 r0 *1 132.8,113.4
X$47 166 163 125 3 pfet_06v0_dn_CDNS_6312644960742
* cell instance $48 r0 *1 146.8,113.4
X$48 168 165 126 3 pfet_06v0_dn_CDNS_6312644960743
* cell instance $49 r0 *1 161.8,113.4
X$49 170 167 127 3 pfet_06v0_dn_CDNS_6312644960744
* cell instance $50 r0 *1 178,113.4
X$50 172 169 128 3 pfet_06v0_dn_CDNS_6312644960745
* cell instance $51 r0 *1 195.6,113.4
X$51 174 171 129 3 pfet_06v0_dn_CDNS_6312644960746
* cell instance $52 r0 *1 214.8,113.4
X$52 176 173 130 3 pfet_06v0_dn_CDNS_6312644960747
* cell instance $53 r0 *1 236,113.4
X$53 178 175 131 3 pfet_06v0_dn_CDNS_6312644960748
* cell instance $54 r0 *1 259.8,113.4
X$54 180 177 132 3 pfet_06v0_dn_CDNS_6312644960749
* cell instance $55 r0 *1 286.4,113.4
X$55 182 179 133 3 pfet_06v0_dn_CDNS_6312644960750
* cell instance $56 r0 *1 316.6,113.4
X$56 184 181 134 3 pfet_06v0_dn_CDNS_6312644960751
* cell instance $57 r0 *1 351,113.4
X$57 186 183 135 3 pfet_06v0_dn_CDNS_6312644960752
* cell instance $58 r0 *1 390.4,113.4
X$58 188 185 136 3 pfet_06v0_dn_CDNS_6312644960753
* cell instance $59 r0 *1 436,113.4
X$59 190 187 137 3 pfet_06v0_dn_CDNS_6312644960754
* cell instance $60 r0 *1 488.8,113.4
X$60 140 189 138 3 pfet_06v0_dn_CDNS_6312644960791
* cell instance $61 r0 *1 2.4,122
X$61 191 192 193 3 pfet_06v0_dn_CDNS_6312644960756
* cell instance $62 r0 *1 12.2,122
X$62 227 225 194 3 pfet_06v0_dn_CDNS_6312644960757
* cell instance $63 r0 *1 21.8,122
X$63 229 226 195 3 pfet_06v0_dn_CDNS_6312644960758
* cell instance $64 r0 *1 31.4,122
X$64 231 228 196 3 pfet_06v0_dn_CDNS_6312644960759
* cell instance $65 r0 *1 41,122
X$65 233 230 197 3 pfet_06v0_dn_CDNS_6312644960760
* cell instance $66 r0 *1 50.8,122
X$66 235 232 198 3 pfet_06v0_dn_CDNS_6312644960761
* cell instance $67 r0 *1 60.4,122
X$67 237 234 199 3 pfet_06v0_dn_CDNS_6312644960762
* cell instance $68 r0 *1 70,122
X$68 239 236 200 3 pfet_06v0_dn_CDNS_6312644960763
* cell instance $69 r0 *1 79.6,122
X$69 241 238 201 3 pfet_06v0_dn_CDNS_6312644960764
* cell instance $70 r0 *1 89.2,122
X$70 243 240 202 3 pfet_06v0_dn_CDNS_6312644960765
* cell instance $71 r0 *1 98.8,122
X$71 245 242 203 3 pfet_06v0_dn_CDNS_6312644960766
* cell instance $72 r0 *1 108.6,122
X$72 247 244 204 3 pfet_06v0_dn_CDNS_6312644960767
* cell instance $73 r0 *1 118.2,122
X$73 249 246 205 3 pfet_06v0_dn_CDNS_6312644960768
* cell instance $74 r0 *1 127.8,122
X$74 251 248 206 3 pfet_06v0_dn_CDNS_6312644960769
* cell instance $75 r0 *1 137.4,122
X$75 253 250 207 3 pfet_06v0_dn_CDNS_6312644960770
* cell instance $76 r0 *1 147,122
X$76 255 252 208 3 pfet_06v0_dn_CDNS_6312644960771
* cell instance $77 r0 *1 156.6,122
X$77 257 254 209 3 pfet_06v0_dn_CDNS_6312644960772
* cell instance $78 r0 *1 166.2,122
X$78 259 256 210 3 pfet_06v0_dn_CDNS_6312644960773
* cell instance $79 r0 *1 176,122
X$79 261 258 211 3 pfet_06v0_dn_CDNS_6312644960774
* cell instance $80 r0 *1 185.6,122
X$80 263 260 212 3 pfet_06v0_dn_CDNS_6312644960775
* cell instance $81 r0 *1 195.2,122
X$81 265 262 213 3 pfet_06v0_dn_CDNS_6312644960776
* cell instance $82 r0 *1 204.8,122
X$82 267 264 214 3 pfet_06v0_dn_CDNS_6312644960777
* cell instance $83 r0 *1 214.4,122
X$83 269 266 215 3 pfet_06v0_dn_CDNS_6312644960778
* cell instance $84 r0 *1 224,122
X$84 271 268 216 3 pfet_06v0_dn_CDNS_6312644960779
* cell instance $85 r0 *1 233.6,122
X$85 270 273 217 3 pfet_06v0_dn_CDNS_6312644960780
* cell instance $86 r0 *1 243.4,122
X$86 272 275 218 3 pfet_06v0_dn_CDNS_6312644960781
* cell instance $87 r0 *1 253,122
X$87 274 277 219 3 pfet_06v0_dn_CDNS_6312644960782
* cell instance $88 r0 *1 262.6,122
X$88 276 279 220 3 pfet_06v0_dn_CDNS_6312644960783
* cell instance $89 r0 *1 272.2,122
X$89 278 281 221 3 pfet_06v0_dn_CDNS_6312644960784
* cell instance $90 r0 *1 281.8,122
X$90 280 283 222 3 pfet_06v0_dn_CDNS_6312644960785
* cell instance $91 r0 *1 291.4,122
X$91 282 285 223 3 pfet_06v0_dn_CDNS_6312644960786
* cell instance $92 r0 *1 301.2,122
X$92 284 287 224 3 pfet_06v0_dn_CDNS_6312644960787
* cell instance $93 r0 *1 310.8,122
X$93 288 286 289 3 pfet_06v0_dn_CDNS_6312644960755
* cell instance $94 r0 *1 2.2,87.6
X$94 90 92 86 3 pfet_06v0_dn_CDNS_6312644960712
* cell instance $95 r0 *1 11.8,61.8
X$95 44 46 39 3 pfet_06v0_dn_CDNS_6312644960713
* cell instance $96 r0 *1 2.2,104.8
X$96 108 107 104 3 pfet_06v0_dn_CDNS_631264496070
* cell instance $97 r0 *1 -34.615,96.2
X$97 100 98 97 3 pfet_06v0_dn_CDNS_631264496070
.ENDS sample_pfet_06v0_dn

* cell M1_NACTIVE_CDNS_631264496070
* pin 
.SUBCKT M1_NACTIVE_CDNS_631264496070 1
.ENDS M1_NACTIVE_CDNS_631264496070

* cell pfet_06v0_dn_CDNS_6312644960791
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960791 1 3 4 6
* device instance $1 r0 *1 25,0.18 pfet_06v0_dn
M$1 3 4 1 6 pfet_06v0_dn L=50U W=0.36U AS=0.1584P AD=0.0936P PS=1.6U PD=0.88U
* device instance $2 r0 *1 75.52,0.18 pfet_06v0_dn
M$2 1 4 3 6 pfet_06v0_dn L=50U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $3 r0 *1 126.04,0.18 pfet_06v0_dn
M$3 3 4 1 6 pfet_06v0_dn L=50U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $4 r0 *1 176.56,0.18 pfet_06v0_dn
M$4 1 4 3 6 pfet_06v0_dn L=50U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $5 r0 *1 227.08,0.18 pfet_06v0_dn
M$5 3 4 1 6 pfet_06v0_dn L=50U W=0.36U AS=0.0936P AD=0.1584P PS=0.88U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960791

* cell pfet_06v0_dn_CDNS_6312644960790
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960790 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.0936P PS=1.6U PD=0.88U
* device instance $2 r0 *1 1.345,0.18 pfet_06v0_dn
M$2 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.1584P PS=0.88U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960790

* cell pfet_06v0_dn_CDNS_6312644960789
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960789 1 4 5 6
* device instance $1 r0 *1 0.275,4.18 pfet_06v0_dn
M$1 5 6 4 1 pfet_06v0_dn L=0.55U W=8.36U AS=3.6784P AD=2.1736P PS=17.6U PD=8.88U
* device instance $2 r0 *1 1.345,4.18 pfet_06v0_dn
M$2 4 6 5 1 pfet_06v0_dn L=0.55U W=8.36U AS=2.1736P AD=2.1736P PS=8.88U PD=8.88U
* device instance $3 r0 *1 2.415,4.18 pfet_06v0_dn
M$3 5 6 4 1 pfet_06v0_dn L=0.55U W=8.36U AS=2.1736P AD=3.6784P PS=8.88U PD=17.6U
.ENDS pfet_06v0_dn_CDNS_6312644960789

* cell pfet_06v0_dn_CDNS_6312644960788
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960788 3 4 5 6
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 5 6 4 3 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960788

* cell pfet_06v0_dn_CDNS_6312644960787
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960787 2 3 4 5
* device instance $1 r0 *1 0.275,42.727 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=85.455U AS=37.6002P AD=37.6002P PS=171.79U
+ PD=171.79U
.ENDS pfet_06v0_dn_CDNS_6312644960787

* cell pfet_06v0_dn_CDNS_6312644960786
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960786 2 3 4 5
* device instance $1 r0 *1 0.275,35.607 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=71.215U AS=31.3346P AD=31.3346P PS=143.31U
+ PD=143.31U
.ENDS pfet_06v0_dn_CDNS_6312644960786

* cell pfet_06v0_dn_CDNS_6312644960785
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960785 2 3 4 5
* device instance $1 r0 *1 0.275,29.672 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=59.345U AS=26.1118P AD=26.1118P PS=119.57U
+ PD=119.57U
.ENDS pfet_06v0_dn_CDNS_6312644960785

* cell pfet_06v0_dn_CDNS_6312644960784
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960784 2 3 4 5
* device instance $1 r0 *1 0.275,24.727 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=49.455U AS=21.7602P AD=21.7602P PS=99.79U
+ PD=99.79U
.ENDS pfet_06v0_dn_CDNS_6312644960784

* cell pfet_06v0_dn_CDNS_6312644960783
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960783 2 3 4 5
* device instance $1 r0 *1 0.275,20.605 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=41.21U AS=18.1324P AD=18.1324P PS=83.3U
+ PD=83.3U
.ENDS pfet_06v0_dn_CDNS_6312644960783

* cell pfet_06v0_dn_CDNS_6312644960782
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960782 2 3 4 5
* device instance $1 r0 *1 0.275,17.172 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=34.345U AS=15.1118P AD=15.1118P PS=69.57U
+ PD=69.57U
.ENDS pfet_06v0_dn_CDNS_6312644960782

* cell pfet_06v0_dn_CDNS_6312644960781
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960781 2 3 4 5
* device instance $1 r0 *1 0.275,14.31 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=28.62U AS=12.5928P AD=12.5928P PS=58.12U
+ PD=58.12U
.ENDS pfet_06v0_dn_CDNS_6312644960781

* cell pfet_06v0_dn_CDNS_6312644960780
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960780 2 3 4 5
* device instance $1 r0 *1 0.275,11.925 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=23.85U AS=10.494P AD=10.494P PS=48.58U
+ PD=48.58U
.ENDS pfet_06v0_dn_CDNS_6312644960780

* cell pfet_06v0_dn_CDNS_6312644960779
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960779 2 3 4 5
* device instance $1 r0 *1 0.275,9.937 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=19.875U AS=8.745P AD=8.745P PS=40.63U
+ PD=40.63U
.ENDS pfet_06v0_dn_CDNS_6312644960779

* cell pfet_06v0_dn_CDNS_6312644960778
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960778 2 3 4 5
* device instance $1 r0 *1 0.275,8.28 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=16.56U AS=7.2864P AD=7.2864P PS=34U PD=34U
.ENDS pfet_06v0_dn_CDNS_6312644960778

* cell pfet_06v0_dn_CDNS_6312644960777
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960777 2 3 4 5
* device instance $1 r0 *1 0.275,6.9 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=13.8U AS=6.072P AD=6.072P PS=28.48U PD=28.48U
.ENDS pfet_06v0_dn_CDNS_6312644960777

* cell pfet_06v0_dn_CDNS_6312644960776
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960776 2 3 4 5
* device instance $1 r0 *1 0.275,5.75 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=11.5U AS=5.06P AD=5.06P PS=23.88U PD=23.88U
.ENDS pfet_06v0_dn_CDNS_6312644960776

* cell pfet_06v0_dn_CDNS_6312644960775
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960775 2 3 4 5
* device instance $1 r0 *1 0.275,4.792 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=9.585U AS=4.2174P AD=4.2174P PS=20.05U
+ PD=20.05U
.ENDS pfet_06v0_dn_CDNS_6312644960775

* cell pfet_06v0_dn_CDNS_6312644960774
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960774 2 3 4 5
* device instance $1 r0 *1 0.275,3.992 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=7.985U AS=3.5134P AD=3.5134P PS=16.85U
+ PD=16.85U
.ENDS pfet_06v0_dn_CDNS_6312644960774

* cell pfet_06v0_dn_CDNS_6312644960773
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960773 2 3 4 5
* device instance $1 r0 *1 0.275,3.327 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=6.655U AS=2.9282P AD=2.9282P PS=14.19U
+ PD=14.19U
.ENDS pfet_06v0_dn_CDNS_6312644960773

* cell pfet_06v0_dn_CDNS_6312644960772
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960772 2 3 4 5
* device instance $1 r0 *1 0.275,2.772 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=5.545U AS=2.4398P AD=2.4398P PS=11.97U
+ PD=11.97U
.ENDS pfet_06v0_dn_CDNS_6312644960772

* cell pfet_06v0_dn_CDNS_6312644960771
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960771 2 3 4 5
* device instance $1 r0 *1 0.275,2.31 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=4.62U AS=2.0328P AD=2.0328P PS=10.12U
+ PD=10.12U
.ENDS pfet_06v0_dn_CDNS_6312644960771

* cell pfet_06v0_dn_CDNS_6312644960770
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960770 2 3 4 5
* device instance $1 r0 *1 0.275,1.925 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=3.85U AS=1.694P AD=1.694P PS=8.58U PD=8.58U
.ENDS pfet_06v0_dn_CDNS_6312644960770

* cell pfet_06v0_dn_CDNS_6312644960769
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960769 2 3 4 5
* device instance $1 r0 *1 0.275,1.605 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=3.21U AS=1.4124P AD=1.4124P PS=7.3U PD=7.3U
.ENDS pfet_06v0_dn_CDNS_6312644960769

* cell pfet_06v0_dn_CDNS_6312644960768
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960768 2 3 4 5
* device instance $1 r0 *1 0.275,1.337 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=2.675U AS=1.177P AD=1.177P PS=6.23U PD=6.23U
.ENDS pfet_06v0_dn_CDNS_6312644960768

* cell pfet_06v0_dn_CDNS_6312644960767
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960767 2 3 4 5
* device instance $1 r0 *1 0.275,1.115 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=2.23U AS=0.9812P AD=0.9812P PS=5.34U PD=5.34U
.ENDS pfet_06v0_dn_CDNS_6312644960767

* cell pfet_06v0_dn_CDNS_6312644960766
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960766 2 3 4 5
* device instance $1 r0 *1 0.275,0.93 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=1.86U AS=0.8184P AD=0.8184P PS=4.6U PD=4.6U
.ENDS pfet_06v0_dn_CDNS_6312644960766

* cell pfet_06v0_dn_CDNS_6312644960765
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960765 2 3 4 5
* device instance $1 r0 *1 0.275,0.775 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=1.55U AS=0.682P AD=0.682P PS=3.98U PD=3.98U
.ENDS pfet_06v0_dn_CDNS_6312644960765

* cell pfet_06v0_dn_CDNS_6312644960764
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960764 2 3 4 5
* device instance $1 r0 *1 0.275,0.645 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=1.29U AS=0.5676P AD=0.5676P PS=3.46U PD=3.46U
.ENDS pfet_06v0_dn_CDNS_6312644960764

* cell pfet_06v0_dn_CDNS_6312644960763
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960763 2 3 4 5
* device instance $1 r0 *1 0.275,0.537 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=1.075U AS=0.473P AD=0.473P PS=3.03U PD=3.03U
.ENDS pfet_06v0_dn_CDNS_6312644960763

* cell pfet_06v0_dn_CDNS_6312644960762
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960762 2 3 4 5
* device instance $1 r0 *1 0.275,0.447 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.895U AS=0.3938P AD=0.3938P PS=2.67U
+ PD=2.67U
.ENDS pfet_06v0_dn_CDNS_6312644960762

* cell pfet_06v0_dn_CDNS_6312644960761
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960761 2 3 4 5
* device instance $1 r0 *1 0.275,0.372 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.745U AS=0.3278P AD=0.3278P PS=2.37U
+ PD=2.37U
.ENDS pfet_06v0_dn_CDNS_6312644960761

* cell pfet_06v0_dn_CDNS_6312644960760
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960760 2 3 4 5
* device instance $1 r0 *1 0.275,0.31 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.62U AS=0.2728P AD=0.2728P PS=2.12U PD=2.12U
.ENDS pfet_06v0_dn_CDNS_6312644960760

* cell pfet_06v0_dn_CDNS_6312644960759
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960759 2 3 4 5
* device instance $1 r0 *1 0.275,0.26 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.52U AS=0.2288P AD=0.2288P PS=1.92U PD=1.92U
.ENDS pfet_06v0_dn_CDNS_6312644960759

* cell pfet_06v0_dn_CDNS_6312644960758
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960758 2 3 4 5
* device instance $1 r0 *1 0.275,0.215 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.43U AS=0.1892P AD=0.1892P PS=1.74U PD=1.74U
.ENDS pfet_06v0_dn_CDNS_6312644960758

* cell pfet_06v0_dn_CDNS_6312644960757
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960757 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960757

* cell pfet_06v0_dn_CDNS_6312644960756
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960756 2 3 4 5
* device instance $1 r0 *1 0.275,0.15 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.3U AS=0.2196P AD=0.2196P PS=2.04U PD=2.04U
.ENDS pfet_06v0_dn_CDNS_6312644960756

* cell pfet_06v0_dn_CDNS_6312644960755
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960755 1 3 4 7
* device instance $1 r0 *1 0.275,50 pfet_06v0_dn
M$1 3 4 1 7 pfet_06v0_dn L=0.55U W=100U AS=44P AD=26P PS=200.88U PD=100.52U
* device instance $2 r0 *1 1.345,50 pfet_06v0_dn
M$2 1 4 3 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $3 r0 *1 2.415,50 pfet_06v0_dn
M$3 3 4 1 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $4 r0 *1 3.485,50 pfet_06v0_dn
M$4 1 4 3 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $5 r0 *1 4.555,50 pfet_06v0_dn
M$5 3 4 1 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $6 r0 *1 5.625,50 pfet_06v0_dn
M$6 1 4 3 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $7 r0 *1 6.695,50 pfet_06v0_dn
M$7 3 4 1 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $8 r0 *1 7.765,50 pfet_06v0_dn
M$8 1 4 3 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $9 r0 *1 8.835,50 pfet_06v0_dn
M$9 3 4 1 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=26P PS=100.52U PD=100.52U
* device instance $10 r0 *1 9.905,50 pfet_06v0_dn
M$10 1 4 3 7 pfet_06v0_dn L=0.55U W=100U AS=26P AD=44P PS=100.52U PD=200.88U
.ENDS pfet_06v0_dn_CDNS_6312644960755

* cell pfet_06v0_dn_CDNS_6312644960754
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960754 2 3 4 5
* device instance $1 r0 *1 21.862,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=43.725U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960754

* cell pfet_06v0_dn_CDNS_6312644960753
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960753 2 3 4 5
* device instance $1 r0 *1 18.217,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=36.435U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960753

* cell pfet_06v0_dn_CDNS_6312644960752
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960752 2 3 4 5
* device instance $1 r0 *1 15.182,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=30.365U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960752

* cell pfet_06v0_dn_CDNS_6312644960751
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960751 2 3 4 5
* device instance $1 r0 *1 12.652,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=25.305U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960751

* cell pfet_06v0_dn_CDNS_6312644960750
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960750 2 3 4 5
* device instance $1 r0 *1 10.542,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=21.085U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960750

* cell pfet_06v0_dn_CDNS_6312644960749
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960749 2 3 4 5
* device instance $1 r0 *1 8.785,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=17.57U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960749

* cell pfet_06v0_dn_CDNS_6312644960748
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960748 2 3 4 5
* device instance $1 r0 *1 7.322,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=14.645U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960748

* cell pfet_06v0_dn_CDNS_6312644960747
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960747 2 3 4 5
* device instance $1 r0 *1 6.1,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=12.2U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960747

* cell pfet_06v0_dn_CDNS_6312644960746
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960746 2 3 4 5
* device instance $1 r0 *1 5.085,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=10.17U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960746

* cell pfet_06v0_dn_CDNS_6312644960745
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960745 2 3 4 5
* device instance $1 r0 *1 4.237,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=8.475U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960745

* cell pfet_06v0_dn_CDNS_6312644960744
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960744 2 3 4 5
* device instance $1 r0 *1 3.53,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=7.06U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960744

* cell pfet_06v0_dn_CDNS_6312644960743
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960743 2 3 4 5
* device instance $1 r0 *1 2.942,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=5.885U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960743

* cell pfet_06v0_dn_CDNS_6312644960742
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960742 2 3 4 5
* device instance $1 r0 *1 2.452,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=4.905U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960742

* cell pfet_06v0_dn_CDNS_6312644960741
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960741 2 3 4 5
* device instance $1 r0 *1 2.042,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=4.085U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960741

* cell pfet_06v0_dn_CDNS_6312644960740
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960740 2 3 4 5
* device instance $1 r0 *1 1.702,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=3.405U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960740

* cell pfet_06v0_dn_CDNS_6312644960739
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960739 2 3 4 5
* device instance $1 r0 *1 1.42,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=2.84U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960739

* cell pfet_06v0_dn_CDNS_6312644960738
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960738 2 3 4 5
* device instance $1 r0 *1 1.182,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=2.365U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960738

* cell pfet_06v0_dn_CDNS_6312644960737
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960737 2 3 4 5
* device instance $1 r0 *1 0.985,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=1.97U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960737

* cell pfet_06v0_dn_CDNS_6312644960736
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960736 2 3 4 5
* device instance $1 r0 *1 0.82,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=1.64U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960736

* cell pfet_06v0_dn_CDNS_6312644960735
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960735 2 3 4 5
* device instance $1 r0 *1 0.685,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=1.37U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960735

* cell pfet_06v0_dn_CDNS_6312644960734
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960734 2 3 4 5
* device instance $1 r0 *1 0.57,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=1.14U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960734

* cell pfet_06v0_dn_CDNS_6312644960733
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960733 2 3 4 5
* device instance $1 r0 *1 0.475,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.95U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960733

* cell pfet_06v0_dn_CDNS_6312644960732
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960732 2 3 4 5
* device instance $1 r0 *1 0.395,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.79U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960732

* cell pfet_06v0_dn_CDNS_6312644960731
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960731 2 3 4 5
* device instance $1 r0 *1 0.33,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.66U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960731

* cell pfet_06v0_dn_CDNS_6312644960730
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960730 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960730

* cell pfet_06v0_dn_CDNS_6312644960729
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960729 1 3 4 8
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.0936P PS=1.6U PD=0.88U
* device instance $2 r0 *1 1.345,0.18 pfet_06v0_dn
M$2 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $3 r0 *1 2.415,0.18 pfet_06v0_dn
M$3 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $4 r0 *1 3.485,0.18 pfet_06v0_dn
M$4 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $5 r0 *1 4.555,0.18 pfet_06v0_dn
M$5 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $6 r0 *1 5.625,0.18 pfet_06v0_dn
M$6 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $7 r0 *1 6.695,0.18 pfet_06v0_dn
M$7 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $8 r0 *1 7.765,0.18 pfet_06v0_dn
M$8 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $9 r0 *1 8.835,0.18 pfet_06v0_dn
M$9 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $10 r0 *1 9.905,0.18 pfet_06v0_dn
M$10 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $11 r0 *1 10.975,0.18 pfet_06v0_dn
M$11 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $12 r0 *1 12.045,0.18 pfet_06v0_dn
M$12 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $13 r0 *1 13.115,0.18 pfet_06v0_dn
M$13 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $14 r0 *1 14.185,0.18 pfet_06v0_dn
M$14 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $15 r0 *1 15.255,0.18 pfet_06v0_dn
M$15 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $16 r0 *1 16.325,0.18 pfet_06v0_dn
M$16 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $17 r0 *1 17.395,0.18 pfet_06v0_dn
M$17 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $18 r0 *1 18.465,0.18 pfet_06v0_dn
M$18 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $19 r0 *1 19.535,0.18 pfet_06v0_dn
M$19 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $20 r0 *1 20.605,0.18 pfet_06v0_dn
M$20 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $21 r0 *1 21.675,0.18 pfet_06v0_dn
M$21 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $22 r0 *1 22.745,0.18 pfet_06v0_dn
M$22 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $23 r0 *1 23.815,0.18 pfet_06v0_dn
M$23 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $24 r0 *1 24.885,0.18 pfet_06v0_dn
M$24 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $25 r0 *1 25.955,0.18 pfet_06v0_dn
M$25 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $26 r0 *1 27.025,0.18 pfet_06v0_dn
M$26 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $27 r0 *1 28.095,0.18 pfet_06v0_dn
M$27 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $28 r0 *1 29.165,0.18 pfet_06v0_dn
M$28 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $29 r0 *1 30.235,0.18 pfet_06v0_dn
M$29 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $30 r0 *1 31.305,0.18 pfet_06v0_dn
M$30 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $31 r0 *1 32.375,0.18 pfet_06v0_dn
M$31 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $32 r0 *1 33.445,0.18 pfet_06v0_dn
M$32 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $33 r0 *1 34.515,0.18 pfet_06v0_dn
M$33 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $34 r0 *1 35.585,0.18 pfet_06v0_dn
M$34 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $35 r0 *1 36.655,0.18 pfet_06v0_dn
M$35 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $36 r0 *1 37.725,0.18 pfet_06v0_dn
M$36 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $37 r0 *1 38.795,0.18 pfet_06v0_dn
M$37 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $38 r0 *1 39.865,0.18 pfet_06v0_dn
M$38 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $39 r0 *1 40.935,0.18 pfet_06v0_dn
M$39 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $40 r0 *1 42.005,0.18 pfet_06v0_dn
M$40 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $41 r0 *1 43.075,0.18 pfet_06v0_dn
M$41 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $42 r0 *1 44.145,0.18 pfet_06v0_dn
M$42 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $43 r0 *1 45.215,0.18 pfet_06v0_dn
M$43 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $44 r0 *1 46.285,0.18 pfet_06v0_dn
M$44 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $45 r0 *1 47.355,0.18 pfet_06v0_dn
M$45 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $46 r0 *1 48.425,0.18 pfet_06v0_dn
M$46 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $47 r0 *1 49.495,0.18 pfet_06v0_dn
M$47 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $48 r0 *1 50.565,0.18 pfet_06v0_dn
M$48 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $49 r0 *1 51.635,0.18 pfet_06v0_dn
M$49 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $50 r0 *1 52.705,0.18 pfet_06v0_dn
M$50 1 4 3 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $51 r0 *1 53.775,0.18 pfet_06v0_dn
M$51 3 4 1 8 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.1584P PS=0.88U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960729

* cell pfet_06v0_dn_CDNS_6312644960728
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960728 2 3 4 5
* device instance $1 r0 *1 0.275,18 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=36U AS=15.84P AD=15.84P PS=72.88U PD=72.88U
.ENDS pfet_06v0_dn_CDNS_6312644960728

* cell pfet_06v0_dn_CDNS_6312644960727
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960727 3 4 5 6
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 5 6 4 3 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960727

* cell pfet_06v0_dn_CDNS_6312644960726
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960726 2 3 4 5
* device instance $1 r0 *1 0.275,0.15 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=0.3U AS=0.2196P AD=0.1548P PS=2.04U PD=1.32U
* device instance $2 r0 *1 1.785,0.15 pfet_06v0_dn
M$2 3 4 2 5 pfet_06v0_dn L=0.55U W=0.3U AS=0.1548P AD=0.1548P PS=1.32U PD=1.32U
* device instance $3 r0 *1 3.295,0.15 pfet_06v0_dn
M$3 2 4 3 5 pfet_06v0_dn L=0.55U W=0.3U AS=0.1548P AD=0.2196P PS=1.32U PD=2.04U
.ENDS pfet_06v0_dn_CDNS_6312644960726

* cell pfet_06v0_dn_CDNS_6312644960725
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960725 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960725

* cell pfet_06v0_dn_CDNS_6312644960724
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960724 1 3 5 9
* device instance $1 r0 *1 0.275,2.68 pfet_06v0_dn
M$1 5 1 3 9 pfet_06v0_dn L=0.55U W=5.36U AS=2.3584P AD=1.3936P PS=11.6U PD=5.88U
* device instance $2 r0 *1 1.345,2.68 pfet_06v0_dn
M$2 3 1 5 9 pfet_06v0_dn L=0.55U W=5.36U AS=1.3936P AD=1.3936P PS=5.88U PD=5.88U
* device instance $3 r0 *1 2.415,2.68 pfet_06v0_dn
M$3 5 1 3 9 pfet_06v0_dn L=0.55U W=5.36U AS=1.3936P AD=2.3584P PS=5.88U PD=11.6U
.ENDS pfet_06v0_dn_CDNS_6312644960724

* cell pfet_06v0_dn_CDNS_6312644960723
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960723 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.432P AD=0.432P PS=3.12U PD=3.12U
.ENDS pfet_06v0_dn_CDNS_6312644960723

* cell pfet_06v0_dn_CDNS_6312644960722
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960722 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.3726P AD=0.3726P PS=2.79U PD=2.79U
.ENDS pfet_06v0_dn_CDNS_6312644960722

* cell pfet_06v0_dn_CDNS_6312644960721
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960721 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.3222P AD=0.3222P PS=2.51U PD=2.51U
.ENDS pfet_06v0_dn_CDNS_6312644960721

* cell pfet_06v0_dn_CDNS_6312644960720
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960720 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.2808P AD=0.2808P PS=2.28U PD=2.28U
.ENDS pfet_06v0_dn_CDNS_6312644960720

* cell pfet_06v0_dn_CDNS_6312644960719
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960719 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.2466P AD=0.2466P PS=2.09U PD=2.09U
.ENDS pfet_06v0_dn_CDNS_6312644960719

* cell pfet_06v0_dn_CDNS_6312644960718
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960718 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.2178P AD=0.2178P PS=1.93U PD=1.93U
.ENDS pfet_06v0_dn_CDNS_6312644960718

* cell pfet_06v0_dn_CDNS_6312644960717
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960717 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1944P AD=0.1944P PS=1.8U PD=1.8U
.ENDS pfet_06v0_dn_CDNS_6312644960717

* cell pfet_06v0_dn_CDNS_6312644960716
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960716 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1746P AD=0.1746P PS=1.69U PD=1.69U
.ENDS pfet_06v0_dn_CDNS_6312644960716

* cell pfet_06v0_dn_CDNS_6312644960715
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960715 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960715

* cell pfet_06v0_dn_CDNS_6312644960714
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960714 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960714

* cell pfet_06v0_dn_CDNS_6312644960713
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960713 2 3 4 5
* device instance $1 r0 *1 0.275,1.68 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=3.36U AS=1.4784P AD=0.8736P PS=7.6U PD=3.88U
* device instance $2 r0 *1 1.345,1.68 pfet_06v0_dn
M$2 3 4 2 5 pfet_06v0_dn L=0.55U W=3.36U AS=0.8736P AD=1.4784P PS=3.88U PD=7.6U
.ENDS pfet_06v0_dn_CDNS_6312644960713

* cell pfet_06v0_dn_CDNS_6312644960712
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960712 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 2 4 3 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.0936P PS=1.6U PD=0.88U
* device instance $2 r0 *1 1.345,0.18 pfet_06v0_dn
M$2 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $3 r0 *1 2.415,0.18 pfet_06v0_dn
M$3 2 4 3 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.1584P PS=0.88U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960712

* cell pfet_06v0_dn_CDNS_6312644960711
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960711 1 3 4 7
* device instance $1 r0 *1 0.275,2.68 pfet_06v0_dn
M$1 3 4 1 7 pfet_06v0_dn L=0.55U W=5.36U AS=6.4856P AD=3.4572P PS=13.14U
+ PD=6.65U
* device instance $2 r0 *1 2.115,2.68 pfet_06v0_dn
M$2 1 4 3 7 pfet_06v0_dn L=0.55U W=5.36U AS=3.4572P AD=3.4572P PS=6.65U PD=6.65U
* device instance $3 r0 *1 3.955,2.68 pfet_06v0_dn
M$3 3 4 1 7 pfet_06v0_dn L=0.55U W=5.36U AS=3.4572P AD=3.4572P PS=6.65U PD=6.65U
* device instance $4 r0 *1 5.795,2.68 pfet_06v0_dn
M$4 1 4 3 7 pfet_06v0_dn L=0.55U W=5.36U AS=3.4572P AD=3.4572P PS=6.65U PD=6.65U
* device instance $5 r0 *1 7.635,2.68 pfet_06v0_dn
M$5 3 4 1 7 pfet_06v0_dn L=0.55U W=5.36U AS=3.4572P AD=6.4856P PS=6.65U
+ PD=13.14U
.ENDS pfet_06v0_dn_CDNS_6312644960711

* cell pfet_06v0_dn_CDNS_6312644960710
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_6312644960710 1 3 4 6
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.0936P PS=1.6U PD=0.88U
* device instance $2 r0 *1 1.345,0.18 pfet_06v0_dn
M$2 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $3 r0 *1 2.415,0.18 pfet_06v0_dn
M$3 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $4 r0 *1 3.485,0.18 pfet_06v0_dn
M$4 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $5 r0 *1 4.555,0.18 pfet_06v0_dn
M$5 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $6 r0 *1 5.625,0.18 pfet_06v0_dn
M$6 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $7 r0 *1 6.695,0.18 pfet_06v0_dn
M$7 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $8 r0 *1 7.765,0.18 pfet_06v0_dn
M$8 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $9 r0 *1 8.835,0.18 pfet_06v0_dn
M$9 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U PD=0.88U
* device instance $10 r0 *1 9.905,0.18 pfet_06v0_dn
M$10 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $11 r0 *1 10.975,0.18 pfet_06v0_dn
M$11 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $12 r0 *1 12.045,0.18 pfet_06v0_dn
M$12 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $13 r0 *1 13.115,0.18 pfet_06v0_dn
M$13 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $14 r0 *1 14.185,0.18 pfet_06v0_dn
M$14 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $15 r0 *1 15.255,0.18 pfet_06v0_dn
M$15 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $16 r0 *1 16.325,0.18 pfet_06v0_dn
M$16 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $17 r0 *1 17.395,0.18 pfet_06v0_dn
M$17 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $18 r0 *1 18.465,0.18 pfet_06v0_dn
M$18 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $19 r0 *1 19.535,0.18 pfet_06v0_dn
M$19 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $20 r0 *1 20.605,0.18 pfet_06v0_dn
M$20 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $21 r0 *1 21.675,0.18 pfet_06v0_dn
M$21 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $22 r0 *1 22.745,0.18 pfet_06v0_dn
M$22 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $23 r0 *1 23.815,0.18 pfet_06v0_dn
M$23 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $24 r0 *1 24.885,0.18 pfet_06v0_dn
M$24 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $25 r0 *1 25.955,0.18 pfet_06v0_dn
M$25 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $26 r0 *1 27.025,0.18 pfet_06v0_dn
M$26 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $27 r0 *1 28.095,0.18 pfet_06v0_dn
M$27 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $28 r0 *1 29.165,0.18 pfet_06v0_dn
M$28 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $29 r0 *1 30.235,0.18 pfet_06v0_dn
M$29 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $30 r0 *1 31.305,0.18 pfet_06v0_dn
M$30 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $31 r0 *1 32.375,0.18 pfet_06v0_dn
M$31 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $32 r0 *1 33.445,0.18 pfet_06v0_dn
M$32 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $33 r0 *1 34.515,0.18 pfet_06v0_dn
M$33 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $34 r0 *1 35.585,0.18 pfet_06v0_dn
M$34 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $35 r0 *1 36.655,0.18 pfet_06v0_dn
M$35 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $36 r0 *1 37.725,0.18 pfet_06v0_dn
M$36 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $37 r0 *1 38.795,0.18 pfet_06v0_dn
M$37 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $38 r0 *1 39.865,0.18 pfet_06v0_dn
M$38 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $39 r0 *1 40.935,0.18 pfet_06v0_dn
M$39 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $40 r0 *1 42.005,0.18 pfet_06v0_dn
M$40 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $41 r0 *1 43.075,0.18 pfet_06v0_dn
M$41 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $42 r0 *1 44.145,0.18 pfet_06v0_dn
M$42 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $43 r0 *1 45.215,0.18 pfet_06v0_dn
M$43 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $44 r0 *1 46.285,0.18 pfet_06v0_dn
M$44 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $45 r0 *1 47.355,0.18 pfet_06v0_dn
M$45 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $46 r0 *1 48.425,0.18 pfet_06v0_dn
M$46 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $47 r0 *1 49.495,0.18 pfet_06v0_dn
M$47 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $48 r0 *1 50.565,0.18 pfet_06v0_dn
M$48 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $49 r0 *1 51.635,0.18 pfet_06v0_dn
M$49 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $50 r0 *1 52.705,0.18 pfet_06v0_dn
M$50 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $51 r0 *1 53.775,0.18 pfet_06v0_dn
M$51 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $52 r0 *1 54.845,0.18 pfet_06v0_dn
M$52 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $53 r0 *1 55.915,0.18 pfet_06v0_dn
M$53 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $54 r0 *1 56.985,0.18 pfet_06v0_dn
M$54 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $55 r0 *1 58.055,0.18 pfet_06v0_dn
M$55 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $56 r0 *1 59.125,0.18 pfet_06v0_dn
M$56 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $57 r0 *1 60.195,0.18 pfet_06v0_dn
M$57 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $58 r0 *1 61.265,0.18 pfet_06v0_dn
M$58 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $59 r0 *1 62.335,0.18 pfet_06v0_dn
M$59 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $60 r0 *1 63.405,0.18 pfet_06v0_dn
M$60 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $61 r0 *1 64.475,0.18 pfet_06v0_dn
M$61 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $62 r0 *1 65.545,0.18 pfet_06v0_dn
M$62 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $63 r0 *1 66.615,0.18 pfet_06v0_dn
M$63 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $64 r0 *1 67.685,0.18 pfet_06v0_dn
M$64 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $65 r0 *1 68.755,0.18 pfet_06v0_dn
M$65 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $66 r0 *1 69.825,0.18 pfet_06v0_dn
M$66 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $67 r0 *1 70.895,0.18 pfet_06v0_dn
M$67 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $68 r0 *1 71.965,0.18 pfet_06v0_dn
M$68 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $69 r0 *1 73.035,0.18 pfet_06v0_dn
M$69 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $70 r0 *1 74.105,0.18 pfet_06v0_dn
M$70 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $71 r0 *1 75.175,0.18 pfet_06v0_dn
M$71 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $72 r0 *1 76.245,0.18 pfet_06v0_dn
M$72 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $73 r0 *1 77.315,0.18 pfet_06v0_dn
M$73 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $74 r0 *1 78.385,0.18 pfet_06v0_dn
M$74 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $75 r0 *1 79.455,0.18 pfet_06v0_dn
M$75 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $76 r0 *1 80.525,0.18 pfet_06v0_dn
M$76 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $77 r0 *1 81.595,0.18 pfet_06v0_dn
M$77 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $78 r0 *1 82.665,0.18 pfet_06v0_dn
M$78 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $79 r0 *1 83.735,0.18 pfet_06v0_dn
M$79 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $80 r0 *1 84.805,0.18 pfet_06v0_dn
M$80 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $81 r0 *1 85.875,0.18 pfet_06v0_dn
M$81 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $82 r0 *1 86.945,0.18 pfet_06v0_dn
M$82 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $83 r0 *1 88.015,0.18 pfet_06v0_dn
M$83 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $84 r0 *1 89.085,0.18 pfet_06v0_dn
M$84 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $85 r0 *1 90.155,0.18 pfet_06v0_dn
M$85 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $86 r0 *1 91.225,0.18 pfet_06v0_dn
M$86 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $87 r0 *1 92.295,0.18 pfet_06v0_dn
M$87 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $88 r0 *1 93.365,0.18 pfet_06v0_dn
M$88 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $89 r0 *1 94.435,0.18 pfet_06v0_dn
M$89 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $90 r0 *1 95.505,0.18 pfet_06v0_dn
M$90 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $91 r0 *1 96.575,0.18 pfet_06v0_dn
M$91 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $92 r0 *1 97.645,0.18 pfet_06v0_dn
M$92 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $93 r0 *1 98.715,0.18 pfet_06v0_dn
M$93 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $94 r0 *1 99.785,0.18 pfet_06v0_dn
M$94 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $95 r0 *1 100.855,0.18 pfet_06v0_dn
M$95 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $96 r0 *1 101.925,0.18 pfet_06v0_dn
M$96 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $97 r0 *1 102.995,0.18 pfet_06v0_dn
M$97 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $98 r0 *1 104.065,0.18 pfet_06v0_dn
M$98 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $99 r0 *1 105.135,0.18 pfet_06v0_dn
M$99 3 4 1 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.0936P PS=0.88U
+ PD=0.88U
* device instance $100 r0 *1 106.205,0.18 pfet_06v0_dn
M$100 1 4 3 6 pfet_06v0_dn L=0.55U W=0.36U AS=0.0936P AD=0.1584P PS=0.88U
+ PD=1.6U
.ENDS pfet_06v0_dn_CDNS_6312644960710

* cell pfet_06v0_dn_CDNS_631264496079
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496079 2 3 4 5
* device instance $1 r0 *1 0.275,9.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=18.36U AS=8.0784P AD=8.0784P PS=37.6U
+ PD=37.6U
.ENDS pfet_06v0_dn_CDNS_631264496079

* cell pfet_06v0_dn_CDNS_631264496078
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496078 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 5 3 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1692P AD=0.1584P PS=1.66U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496078

* cell pfet_06v0_dn_CDNS_631264496077
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496077 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 5 3 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496077

* cell pfet_06v0_dn_CDNS_631264496076
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496076 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 5 3 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496076

* cell pfet_06v0_dn_CDNS_631264496075
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496075 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 5 3 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496075

* cell pfet_06v0_dn_CDNS_631264496074
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496074 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 5 3 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496074

* cell pfet_06v0_dn_CDNS_631264496073
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496073 1 4 5 6
* device instance $1 r0 *1 0.275,1.68 pfet_06v0_dn
M$1 5 6 4 1 pfet_06v0_dn L=0.55U W=3.36U AS=1.4784P AD=0.8736P PS=7.6U PD=3.88U
* device instance $2 r0 *1 1.345,1.68 pfet_06v0_dn
M$2 4 6 5 1 pfet_06v0_dn L=0.55U W=3.36U AS=0.8736P AD=0.8736P PS=3.88U PD=3.88U
* device instance $3 r0 *1 2.415,1.68 pfet_06v0_dn
M$3 5 6 4 1 pfet_06v0_dn L=0.55U W=3.36U AS=0.8736P AD=1.4784P PS=3.88U PD=7.6U
.ENDS pfet_06v0_dn_CDNS_631264496073

* cell pfet_06v0_dn_CDNS_631264496072
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496072 2 4 5 6
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 4 6 5 2 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496072

* cell pfet_06v0_dn_CDNS_631264496071
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496071 3 4 5 6
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 5 6 4 3 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496071

* cell pfet_06v0_dn_CDNS_631264496070
* pin 
* pin 
* pin 
* pin 
.SUBCKT pfet_06v0_dn_CDNS_631264496070 2 3 4 5
* device instance $1 r0 *1 0.275,0.18 pfet_06v0_dn
M$1 3 4 2 5 pfet_06v0_dn L=0.55U W=0.36U AS=0.1584P AD=0.1584P PS=1.6U PD=1.6U
.ENDS pfet_06v0_dn_CDNS_631264496070
